module add2b(
    input [15:0]a,b,
    output [15:0]y
    );
    
    assign y = a+b;
    
endmodule
